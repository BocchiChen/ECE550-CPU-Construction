module RCA_32bit(a,b,cin,sum);
   input [31:0] a, b;
   input cin;
   //output cout;
   output [31:0] sum;
   wire w1,w2,w3,w4,w5,w6,w7,w8,w9,w10,w11,w12,w13,w14,w15,w16,w17,w18,w19,w20,w21,w22,w23,w24,w25,w26,w27,w28,w29,w30,w31;
	
   full_adder f1(a[0], b[0], cin, sum[0], w1);
   full_adder f2(a[1], b[1], w1, sum[1], w2);
   full_adder f3(a[2], b[2], w2, sum[2], w3);
   full_adder f4(a[3], b[3], w3, sum[3], w4);
   full_adder f5(a[4], b[4], w4, sum[4], w5);
   full_adder f6(a[5], b[5], w5, sum[5], w6);
   full_adder f7(a[6], b[6], w6, sum[6], w7);
   full_adder f8(a[7], b[7], w7, sum[7], w8);
	full_adder f9(a[8], b[8], w8, sum[8], w9);
	full_adder f10(a[9], b[9], w9, sum[9], w10);
	full_adder f11(a[10], b[10], w10, sum[10], w11);
	full_adder f12(a[11], b[11], w11, sum[11], w12);
	full_adder f13(a[12], b[12], w12, sum[12], w13);
	full_adder f14(a[13], b[13], w13, sum[13], w14);
	full_adder f15(a[14], b[14], w14, sum[14], w15);
	full_adder f16(a[15], b[15], w15, sum[15], w16);
	full_adder f17(a[16], b[16], w16, sum[16], w17);
	full_adder f18(a[17], b[17], w17, sum[17], w18);
	full_adder f19(a[18], b[18], w18, sum[18], w19);
	full_adder f20(a[19], b[19], w19, sum[19], w20);
	full_adder f21(a[20], b[20], w20, sum[20], w21);
	full_adder f22(a[21], b[21], w21, sum[21], w22);
	full_adder f23(a[22], b[22], w22, sum[22], w23);
	full_adder f24(a[23], b[23], w23, sum[23], w24);
	full_adder f25(a[24], b[24], w24, sum[24], w25);
	full_adder f26(a[25], b[25], w25, sum[25], w26);
	full_adder f27(a[26], b[26], w26, sum[26], w27);
	full_adder f28(a[27], b[27], w27, sum[27], w28);
	full_adder f29(a[28], b[28], w28, sum[28], w29);
	full_adder f30(a[29], b[29], w29, sum[29], w30);
	full_adder f31(a[30], b[30], w30, sum[30], w31);
	full_adder f32(a[31], b[31], w31, sum[31], cout);
	
endmodule
